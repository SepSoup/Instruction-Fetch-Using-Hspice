*CMOS----SepehrBazmi--------------------------------------------------------------------
.include model.sp

.GLOBAL VDD
VDD VDD 0 1.1
.GLOBAL CLK
VCLK CLK 0 0 PULSE(1.1 0 5p 0.001N 0.001N 100N 200N)


XPC D0 D1 D2 D3 Q0 Q1 Q2 Q3 PC
XALU Q0 Q1 Q2 Q3 D0 D1 D2 D3 ALU
XIM Q0 Q1 Q2 Q3 O31 O30 O29 O28 O27 O26 O25 O24 O23 O22 O21 O20 O19 O18 O17 O16 O15 O14 O13 O12 O11 O10 O9 O8 O7 O6 O5 O4 O3 O2 O1 O0 IM




.TRAN 10P 9U



*---INSTRUCTION-MEMORY---------------------------------------------------------------------------------

.SUBCKT IM IN1 IN2 IN3 IN4 OUT1 OUT2 OUT3 OUT4 OUT5 OUT6 OUT7 OUT8 OUT9 OUT10 OUT11 OUT12 OUT13 OUT14 OUT15 OUT16 OUT17 OUT18 OUT19 OUT20 OUT21 OUT22 OUT23 OUT24 OUT25 OUT26 OUT27 OUT28 OUT29 OUT30 OUT31 OUT32


RC1 VDD C1 100k
RC2 VDD C2 100k
RC3 VDD C3 100k
RC4 VDD C4 100k
RC5 VDD C5 100k
RC6 VDD C6 100k
RC7 VDD C7 100k
RC8 VDD C8 100k
RC9 VDD C9 100k
RC10 VDD C10 100k
RC11 VDD C11 100k
RC12 VDD C12 100k
RC13 VDD C13 100k
RC14 VDD C14 100k
RC15 VDD C15 100k
RC16 VDD C16 100k
RC17 VDD C17 100k
RC18 VDD C18 100k
RC19 VDD C19 100k
RC20 VDD C20 100k
RC21 VDD C21 100k
RC22 VDD C22 100k
RC23 VDD C23 100k
RC24 VDD C24 100k
RC25 VDD C25 100k
RC26 VDD C26 100k
RC27 VDD C27 100k
RC28 VDD C28 100k
RC29 VDD C29 100k
RC30 VDD C30 100k
RC31 VDD C31 100k
RC32 VDD C32 100k

XDEC416 IN1 IN2 IN3 IN4 R1 R2 R3 R4 R5 R6 R7 R8 R9 R10 R11 R12 R13 R14 R15 R16 DEC416


*-------------------------------
MN1 C32 R1 0 0 NMOS L=32N W=1U
MN2 C31 R1 0 0 NMOS L=32N W=1U
*MN3 C30 R1 0 0 NMOS L=32N W=1U
MN4 C29 R1 0 0 NMOS L=32N W=1U
MN5 C28 R1 0 0 NMOS L=32N W=1U
MN6 C27 R1 0 0 NMOS L=32N W=1U
MN7 C26 R1 0 0 NMOS L=32N W=1U
MN8 C25 R1 0 0 NMOS L=32N W=1U
MN9 C24 R1 0 0 NMOS L=32N W=1U
MN10 C23 R1 0 0 NMOS L=32N W=1U
MN11 C22 R1 0 0 NMOS L=32N W=1U
MN12 C21 R1 0 0 NMOS L=32N W=1U
MN13 C20 R1 0 0 NMOS L=32N W=1U
MN14 C19 R1 0 0 NMOS L=32N W=1U
*MN15 C18 R1 0 0 NMOS L=32N W=1U
*MN16 C17 R1 0 0 NMOS L=32N W=1U
MN17 C16 R1 0 0 NMOS L=32N W=1U
MN18 C15 R1 0 0 NMOS L=32N W=1U
MN19 C14 R1 0 0 NMOS L=32N W=1U
MN20 C13 R1 0 0 NMOS L=32N W=1U
MN21 C12 R1 0 0 NMOS L=32N W=1U
MN22 C11 R1 0 0 NMOS L=32N W=1U
MN23 C10 R1 0 0 NMOS L=32N W=1U
MN24 C9 R1 0 0 NMOS L=32N W=1U
MN25 C8 R1 0 0 NMOS L=32N W=1U
MN26 C7 R1 0 0 NMOS L=32N W=1U
MN27 C6 R1 0 0 NMOS L=32N W=1U
MN28 C5 R1 0 0 NMOS L=32N W=1U
*MN29 C4 R1 0 0 NMOS L=32N W=1U
MN30 C3 R1 0 0 NMOS L=32N W=1U
MN31 C2 R1 0 0 NMOS L=32N W=1U
MN32 C1 R1 0 0 NMOS L=32N W=1U
*-------------------------------
MN33 C32 R2 0 0 NMOS L=32N W=1U
MN34 C31 R2 0 0 NMOS L=32N W=1U
*MN35 C30 R2 0 0 NMOS L=32N W=1U
MN36 C29 R2 0 0 NMOS L=32N W=1U
MN37 C28 R2 0 0 NMOS L=32N W=1U
MN38 C27 R2 0 0 NMOS L=32N W=1U
MN39 C26 R2 0 0 NMOS L=32N W=1U
MN40 C25 R2 0 0 NMOS L=32N W=1U
MN41 C24 R2 0 0 NMOS L=32N W=1U
MN42 C23 R2 0 0 NMOS L=32N W=1U
MN43 C22 R2 0 0 NMOS L=32N W=1U
MN44 C21 R2 0 0 NMOS L=32N W=1U
MN45 C20 R2 0 0 NMOS L=32N W=1U
*MN46 C19 R2 0 0 NMOS L=32N W=1U
MN47 C18 R2 0 0 NMOS L=32N W=1U
MN48 C17 R2 0 0 NMOS L=32N W=1U
MN49 C16 R2 0 0 NMOS L=32N W=1U
MN50 C15 R2 0 0 NMOS L=32N W=1U
MN51 C14 R2 0 0 NMOS L=32N W=1U
MN52 C13 R2 0 0 NMOS L=32N W=1U
MN53 C12 R2 0 0 NMOS L=32N W=1U
MN54 C11 R2 0 0 NMOS L=32N W=1U
MN55 C10 R2 0 0 NMOS L=32N W=1U
MN56 C9 R2 0 0 NMOS L=32N W=1U
MN57 C8 R2 0 0 NMOS L=32N W=1U
MN58 C7 R2 0 0 NMOS L=32N W=1U
MN59 C6 R2 0 0 NMOS L=32N W=1U
MN60 C5 R2 0 0 NMOS L=32N W=1U
MN61 C4 R2 0 0 NMOS L=32N W=1U
MN62 C3 R2 0 0 NMOS L=32N W=1U
MN63 C2 R2 0 0 NMOS L=32N W=1U
*MN64 C1 R2 0 0 NMOS L=32N W=1U
*-------------------------------
MN65 C32 R3 0 0 NMOS L=32N W=1U
MN66 C31 R3 0 0 NMOS L=32N W=1U
*MN67 C30 R3 0 0 NMOS L=32N W=1U
MN68 C29 R3 0 0 NMOS L=32N W=1U
MN69 C28 R3 0 0 NMOS L=32N W=1U
MN70 C27 R3 0 0 NMOS L=32N W=1U
MN71 C26 R3 0 0 NMOS L=32N W=1U
MN72 C25 R3 0 0 NMOS L=32N W=1U
MN73 C24 R3 0 0 NMOS L=32N W=1U
MN74 C23 R3 0 0 NMOS L=32N W=1U
MN75 C22 R3 0 0 NMOS L=32N W=1U
MN76 C21 R3 0 0 NMOS L=32N W=1U
MN77 C20 R3 0 0 NMOS L=32N W=1U
*MN78 C19 R3 0 0 NMOS L=32N W=1U
MN79 C18 R3 0 0 NMOS L=32N W=1U
*MN80 C17 R3 0 0 NMOS L=32N W=1U
*MN81 C16 R3 0 0 NMOS L=32N W=1U
*MN82 C15 R3 0 0 NMOS L=32N W=1U
*MN83 C14 R3 0 0 NMOS L=32N W=1U
*MN84 C13 R3 0 0 NMOS L=32N W=1U
*MN85 C12 R3 0 0 NMOS L=32N W=1U
*MN86 C11 R3 0 0 NMOS L=32N W=1U
*MN87 C10 R3 0 0 NMOS L=32N W=1U
*MN88 C9 R3 0 0 NMOS L=32N W=1U
*MN89 C8 R3 0 0 NMOS L=32N W=1U
*MN90 C7 R3 0 0 NMOS L=32N W=1U
*MN91 C6 R3 0 0 NMOS L=32N W=1U
*MN92 C5 R3 0 0 NMOS L=32N W=1U
*MN93 C4 R3 0 0 NMOS L=32N W=1U
*MN94 C3 R3 0 0 NMOS L=32N W=1U
*MN95 C2 R3 0 0 NMOS L=32N W=1U
*MN96 C1 R3 0 0 NMOS L=32N W=1U
*-------------------------------
MN97 C32 R4 0 0 NMOS L=32N W=1U
MN98 C31 R4 0 0 NMOS L=32N W=1U
MN99 C30 R4 0 0 NMOS L=32N W=1U
*MN100 C29 R4 0 0 NMOS L=32N W=1U
MN101 C28 R4 0 0 NMOS L=32N W=1U
MN102 C27 R4 0 0 NMOS L=32N W=1U
MN103 C26 R4 0 0 NMOS L=32N W=1U
MN104 C25 R4 0 0 NMOS L=32N W=1U
MN105 C24 R4 0 0 NMOS L=32N W=1U
*MN106 C23 R4 0 0 NMOS L=32N W=1U
*MN107 C22 R4 0 0 NMOS L=32N W=1U
MN108 C21 R4 0 0 NMOS L=32N W=1U
MN109 C20 R4 0 0 NMOS L=32N W=1U
MN110 C19 R4 0 0 NMOS L=32N W=1U
MN111 C18 R4 0 0 NMOS L=32N W=1U
MN112 C17 R4 0 0 NMOS L=32N W=1U
MN113 C16 R4 0 0 NMOS L=32N W=1U
MN114 C15 R4 0 0 NMOS L=32N W=1U
MN115 C14 R4 0 0 NMOS L=32N W=1U
MN116 C13 R4 0 0 NMOS L=32N W=1U
MN117 C12 R4 0 0 NMOS L=32N W=1U
MN118 C11 R4 0 0 NMOS L=32N W=1U
MN119 C10 R4 0 0 NMOS L=32N W=1U
MN120 C9 R4 0 0 NMOS L=32N W=1U
MN121 C8 R4 0 0 NMOS L=32N W=1U
MN122 C7 R4 0 0 NMOS L=32N W=1U
MN123 C6 R4 0 0 NMOS L=32N W=1U
MN124 C5 R4 0 0 NMOS L=32N W=1U
MN125 C4 R4 0 0 NMOS L=32N W=1U
*MN126 C3 R4 0 0 NMOS L=32N W=1U
MN127 C2 R4 0 0 NMOS L=32N W=1U
MN128 C1 R4 0 0 NMOS L=32N W=1U
*-------------------------------
MN129 C32 R5 0 0 NMOS L=32N W=1U
MN130 C31 R5 0 0 NMOS L=32N W=1U
MN131 C30 R5 0 0 NMOS L=32N W=1U
MN132 C29 R5 0 0 NMOS L=32N W=1U
MN133 C28 R5 0 0 NMOS L=32N W=1U
MN134 C27 R5 0 0 NMOS L=32N W=1U
MN135 C26 R5 0 0 NMOS L=32N W=1U
MN136 C25 R5 0 0 NMOS L=32N W=1U
*MN137 C24 R5 0 0 NMOS L=32N W=1U
MN138 C23 R5 0 0 NMOS L=32N W=1U
MN139 C22 R5 0 0 NMOS L=32N W=1U
MN140 C21 R5 0 0 NMOS L=32N W=1U
MN141 C20 R5 0 0 NMOS L=32N W=1U
*MN142 C19 R5 0 0 NMOS L=32N W=1U
MN143 C18 R5 0 0 NMOS L=32N W=1U
*MN144 C17 R5 0 0 NMOS L=32N W=1U
MN145 C16 R5 0 0 NMOS L=32N W=1U
MN146 C15 R5 0 0 NMOS L=32N W=1U
*MN147 C14 R5 0 0 NMOS L=32N W=1U
MN148 C13 R5 0 0 NMOS L=32N W=1U
MN149 C12 R5 0 0 NMOS L=32N W=1U
MN150 C11 R5 0 0 NMOS L=32N W=1U
MN151 C10 R5 0 0 NMOS L=32N W=1U
MN152 C9 R5 0 0 NMOS L=32N W=1U
MN153 C8 R5 0 0 NMOS L=32N W=1U
MN154 C7 R5 0 0 NMOS L=32N W=1U
*MN155 C6 R5 0 0 NMOS L=32N W=1U
MN156 C5 R5 0 0 NMOS L=32N W=1U
MN157 C4 R5 0 0 NMOS L=32N W=1U
MN158 C3 R5 0 0 NMOS L=32N W=1U
MN159 C2 R5 0 0 NMOS L=32N W=1U
MN160 C1 R5 0 0 NMOS L=32N W=1U
*-------------------------------
MN161 C32 R6 0 0 NMOS L=32N W=1U
MN162 C31 R6 0 0 NMOS L=32N W=1U
MN163 C30 R6 0 0 NMOS L=32N W=1U
MN164 C29 R6 0 0 NMOS L=32N W=1U
MN165 C28 R6 0 0 NMOS L=32N W=1U
MN166 C27 R6 0 0 NMOS L=32N W=1U
MN167 C26 R6 0 0 NMOS L=32N W=1U
MN168 C25 R6 0 0 NMOS L=32N W=1U
*MN169 C24 R6 0 0 NMOS L=32N W=1U
MN170 C23 R6 0 0 NMOS L=32N W=1U
MN171 C22 R6 0 0 NMOS L=32N W=1U
MN172 C21 R6 0 0 NMOS L=32N W=1U
MN173 C20 R6 0 0 NMOS L=32N W=1U
*MN174 C19 R6 0 0 NMOS L=32N W=1U
MN175 C18 R6 0 0 NMOS L=32N W=1U
*MN176 C17 R6 0 0 NMOS L=32N W=1U
MN177 C16 R6 0 0 NMOS L=32N W=1U
MN178 C15 R6 0 0 NMOS L=32N W=1U
*MN179 C14 R6 0 0 NMOS L=32N W=1U
MN180 C13 R6 0 0 NMOS L=32N W=1U
*MN181 C12 R6 0 0 NMOS L=32N W=1U
MN182 C11 R6 0 0 NMOS L=32N W=1U
MN183 C10 R6 0 0 NMOS L=32N W=1U
MN184 C9 R6 0 0 NMOS L=32N W=1U
MN185 C8 R6 0 0 NMOS L=32N W=1U
MN186 C7 R6 0 0 NMOS L=32N W=1U
*MN187 C6 R6 0 0 NMOS L=32N W=1U
MN188 C5 R6 0 0 NMOS L=32N W=1U
MN189 C4 R6 0 0 NMOS L=32N W=1U
MN190 C3 R6 0 0 NMOS L=32N W=1U
*MN191 C2 R6 0 0 NMOS L=32N W=1U
MN192 C1 R6 0 0 NMOS L=32N W=1U
*-------------------------------
MN193 C32 R7 0 0 NMOS L=32N W=1U
MN194 C31 R7 0 0 NMOS L=32N W=1U
*MN195 C30 R7 0 0 NMOS L=32N W=1U
MN196 C29 R7 0 0 NMOS L=32N W=1U
MN197 C28 R7 0 0 NMOS L=32N W=1U
MN198 C27 R7 0 0 NMOS L=32N W=1U
MN199 C26 R7 0 0 NMOS L=32N W=1U
MN200 C25 R7 0 0 NMOS L=32N W=1U
MN201 C24 R7 0 0 NMOS L=32N W=1U
*MN202 C23 R7 0 0 NMOS L=32N W=1U
*MN203 C22 R7 0 0 NMOS L=32N W=1U
MN204 C21 R7 0 0 NMOS L=32N W=1U
MN205 C20 R7 0 0 NMOS L=32N W=1U
MN206 C19 R7 0 0 NMOS L=32N W=1U
*MN207 C18 R7 0 0 NMOS L=32N W=1U
*MN208 C17 R7 0 0 NMOS L=32N W=1U
*MN209 C16 R7 0 0 NMOS L=32N W=1U
*MN210 C15 R7 0 0 NMOS L=32N W=1U
*MN211 C14 R7 0 0 NMOS L=32N W=1U
*MN212 C13 R7 0 0 NMOS L=32N W=1U
*MN213 C12 R7 0 0 NMOS L=32N W=1U
*MN214 C11 R7 0 0 NMOS L=32N W=1U
*MN215 C10 R7 0 0 NMOS L=32N W=1U
*MN216 C9 R7 0 0 NMOS L=32N W=1U
*MN217 C8 R7 0 0 NMOS L=32N W=1U
*MN218 C7 R7 0 0 NMOS L=32N W=1U
*MN219 C6 R7 0 0 NMOS L=32N W=1U
*MN220 C5 R7 0 0 NMOS L=32N W=1U
*MN221 C4 R7 0 0 NMOS L=32N W=1U
*MN222 C3 R7 0 0 NMOS L=32N W=1U
*MN223 C2 R7 0 0 NMOS L=32N W=1U
*MN224 C1 R7 0 0 NMOS L=32N W=1U
*-------------------------------
MN225 C32 R8 0 0 NMOS L=32N W=1U
MN226 C31 R8 0 0 NMOS L=32N W=1U
MN227 C30 R8 0 0 NMOS L=32N W=1U
MN228 C29 R8 0 0 NMOS L=32N W=1U
*MN229 C28 R8 0 0 NMOS L=32N W=1U
MN230 C27 R8 0 0 NMOS L=32N W=1U
MN231 C26 R8 0 0 NMOS L=32N W=1U
MN232 C25 R8 0 0 NMOS L=32N W=1U
MN233 C24 R8 0 0 NMOS L=32N W=1U
MN234 C23 R8 0 0 NMOS L=32N W=1U
MN235 C22 R8 0 0 NMOS L=32N W=1U
MN236 C21 R8 0 0 NMOS L=32N W=1U
MN237 C20 R8 0 0 NMOS L=32N W=1U
MN238 C19 R8 0 0 NMOS L=32N W=1U
MN239 C18 R8 0 0 NMOS L=32N W=1U
MN240 C17 R8 0 0 NMOS L=32N W=1U
MN241 C16 R8 0 0 NMOS L=32N W=1U
MN242 C15 R8 0 0 NMOS L=32N W=1U
MN243 C14 R8 0 0 NMOS L=32N W=1U
MN244 C13 R8 0 0 NMOS L=32N W=1U
MN245 C12 R8 0 0 NMOS L=32N W=1U
MN246 C11 R8 0 0 NMOS L=32N W=1U
MN247 C10 R8 0 0 NMOS L=32N W=1U
MN248 C9 R8 0 0 NMOS L=32N W=1U
MN249 C8 R8 0 0 NMOS L=32N W=1U
MN250 C7 R8 0 0 NMOS L=32N W=1U
MN251 C6 R8 0 0 NMOS L=32N W=1U
MN252 C5 R8 0 0 NMOS L=32N W=1U
MN253 C4 R8 0 0 NMOS L=32N W=1U
MN254 C3 R8 0 0 NMOS L=32N W=1U
*MN255 C2 R8 0 0 NMOS L=32N W=1U
*MN256 C1 R8 0 0 NMOS L=32N W=1U
*-------------------------------
*MN257 C32 R9 0 0 NMOS L=32N W=1U
MN258 C31 R9 0 0 NMOS L=32N W=1U
*MN259 C30 R9 0 0 NMOS L=32N W=1U
MN260 C29 R9 0 0 NMOS L=32N W=1U
MN261 C28 R9 0 0 NMOS L=32N W=1U
MN262 C27 R9 0 0 NMOS L=32N W=1U
MN263 C26 R9 0 0 NMOS L=32N W=1U
MN264 C25 R9 0 0 NMOS L=32N W=1U
MN265 C24 R9 0 0 NMOS L=32N W=1U
MN266 C23 R9 0 0 NMOS L=32N W=1U
MN267 C22 R9 0 0 NMOS L=32N W=1U
MN268 C21 R9 0 0 NMOS L=32N W=1U
MN269 C20 R9 0 0 NMOS L=32N W=1U
*MN270 C19 R9 0 0 NMOS L=32N W=1U
MN271 C18 R9 0 0 NMOS L=32N W=1U
MN272 C17 R9 0 0 NMOS L=32N W=1U
MN273 C16 R9 0 0 NMOS L=32N W=1U
MN274 C15 R9 0 0 NMOS L=32N W=1U
MN275 C14 R9 0 0 NMOS L=32N W=1U
MN276 C13 R9 0 0 NMOS L=32N W=1U
MN277 C12 R9 0 0 NMOS L=32N W=1U
MN278 C11 R9 0 0 NMOS L=32N W=1U
MN279 C10 R9 0 0 NMOS L=32N W=1U
MN280 C9 R9 0 0 NMOS L=32N W=1U
*MN281 C8 R9 0 0 NMOS L=32N W=1U
*MN282 C7 R9 0 0 NMOS L=32N W=1U
*MN283 C6 R9 0 0 NMOS L=32N W=1U
*MN284 C5 R9 0 0 NMOS L=32N W=1U
*MN285 C4 R9 0 0 NMOS L=32N W=1U
*MN286 C3 R9 0 0 NMOS L=32N W=1U
*MN287 C2 R9 0 0 NMOS L=32N W=1U
*MN288 C1 R9 0 0 NMOS L=32N W=1U




XBUFFER1 C1 OUT1 BUFFER
XBUFFER2 C2 OUT2 BUFFER
XBUFFER3 C3 OUT3 BUFFER
XBUFFER4 C4 OUT4 BUFFER
XBUFFER5 C5 OUT5 BUFFER
XBUFFER6 C6 OUT6 BUFFER
XBUFFER7 C7 OUT7 BUFFER
XBUFFER8 C8 OUT8 BUFFER
XBUFFER9 C9 OUT9 BUFFER
XBUFFER10 C10 OUT10 BUFFER
XBUFFER11 C11 OUT11 BUFFER
XBUFFER12 C12 OUT12 BUFFER
XBUFFER13 C13 OUT13 BUFFER
XBUFFER14 C14 OUT14 BUFFER
XBUFFER15 C15 OUT15 BUFFER
XBUFFER16 C16 OUT16 BUFFER
XBUFFER17 C17 OUT17 BUFFER
XBUFFER18 C18 OUT18 BUFFER
XBUFFER19 C19 OUT19 BUFFER
XBUFFER20 C20 OUT20 BUFFER
XBUFFER21 C21 OUT21 BUFFER
XBUFFER22 C22 OUT22 BUFFER
XBUFFER23 C23 OUT23 BUFFER
XBUFFER24 C24 OUT24 BUFFER
XBUFFER25 C25 OUT25 BUFFER
XBUFFER26 C26 OUT26 BUFFER
XBUFFER27 C27 OUT27 BUFFER
XBUFFER28 C28 OUT28 BUFFER
XBUFFER29 C29 OUT29 BUFFER
XBUFFER30 C30 OUT30 BUFFER
XBUFFER31 C31 OUT31 BUFFER
XBUFFER32 C32 OUT32 BUFFER


.ENDS IM

*---NOT---------------------------------------------------------------------------------

.SUBCKT NOT IN OUT 

MP OUT IN VDD VDD PMOS L=32N W=2U
MN OUT IN 0 0 NMOS L=32N W=1U

.ENDS NOT

*---BUFFER---------------------------------------------------------------------------------

.SUBCKT BUFFER IN OUT 

XNOT1 IN NOTIN NOT
XNOT2 NOTIN OUT NOT

.ENDS BUFFER

*---NAND--------------------------------------------------------------------------------

.SUBCKT NAND INA INB OUT 

MP1 OUT INA VDD VDD PMOS L=32N W=2U
MP2 OUT INB VDD VDD PMOS L=32N W=2U

MN1 OUT INA SADB 0 NMOS L=32N W=2U
MN2 SADB INB 0 0 NMOS L=32N W=2U

.ENDS NAND

*---AND---------------------------------------------------------------------------------

.SUBCKT AND INA INB OUT 

XNAND INA INB NANDAB NAND
XNOT NANDAB OUT NOT

.ENDS AND

*---AND3---------------------------------------------------------------------------------

.SUBCKT AND3 INA INB E OUT 

MP1 OUT1 INA VDD VDD PMOS L=32N W=2U
MP2 OUT1 INB VDD VDD PMOS L=32N W=2U
MP3 OUT1 E VDD VDD PMOS L=32N W=2U


MN1 OUT1 INA SMN1 0 NMOS L=32N W=6U
MN2 SMN1 INB SMN2 0 NMOS L=32N W=6U
MN3 SMN2 E 0 0 NMOS L=32N W=6U


XNOT OUT1 OUT NOT


.ENDS AND3


*---AND4---------------------------------------------------------------------------------

.SUBCKT AND4 INA INB INC IND OUT 

MP1 OUT1 INA VDD VDD PMOS L=32N W=2U
MP2 OUT1 INB VDD VDD PMOS L=32N W=2U
MP3 OUT1 INC VDD VDD PMOS L=32N W=2U
MP4 OUT1 IND VDD VDD PMOS L=32N W=2U

MN1 OUT1 INA SMN1 0 NMOS L=32N W=4U
MN2 SMN1 INB SMN2 0 NMOS L=32N W=4U
MN3 SMN2 INC SMN3 0 NMOS L=32N W=4U
MN4 SMN3 IND 0 0 NMOS L=32N W=4U


XNOT OUT1 OUT NOT


.ENDS AND4

*---NOR--------------------------------------------------------------------------------

.SUBCKT NOR INA INB OUT 

MP1 OUT INA SMP1 VDD PMOS L=32N W=2U
MP2 SMP1 INB VDD VDD PMOS L=32N W=2U

MN1 OUT INA 0 0 NMOS L=32N W=2U
MN2 OUT INB 0 0 NMOS L=32N W=2U

.ENDS NOR

*---OR--------------------------------------------------------------------------------

.SUBCKT OR INA INB OUT 

XNOR INA INB NORAB NOR
XNOT NORAB OUT NOT

.ENDS OR


*---XOR--------------------------------------------------------------------------------

.SUBCKT XOR INA INB OUT 

XNOT1 INA NOTA NOT
XNOT2 INB NOTB NOT

XAND1 INA NOTB OUTAND1 AND
XAND2 NOTA INB OUTAND2 AND

XOR OUTAND1 OUTAND2 OUT OR

.ENDS XOR


*---DECODER416--------------------------------------------------------------------------------

.SUBCKT DEC416 IN1 IN2 IN3 IN4 O0 O1 O2 O3 O4 O5 O6 O7 O8 O9 O10 O11 O12 O13 O14 O15

XNOT1 IN1 NOT1 NOT
XNOT2 IN2 NOT2 NOT
XNOT3 IN3 NOT3 NOT
XNOT4 IN4 NOT4 NOT

XAND1 NOT1 NOT2 NOT3 NOT4 O0 AND4
XAND2 IN1 NOT2 NOT3 NOT4 O1 AND4
XAND3 NOT1 IN2 NOT3 NOT4 O2 AND4
XAND4 IN1 IN2 NOT3 NOT4 O3 AND4
XAND5 NOT1 NOT2 IN3 NOT4 O4 AND4
XAND6 IN1 NOT2 IN3 NOT4 O5 AND4
XAND7 NOT1 IN2 IN3 NOT4 O6 AND4
XAND8 IN1 IN2 IN3 NOT4 O7 AND4

XAND9 NOT1 NOT2 NOT3 IN4 O8 AND4
XAND10 IN1 NOT2 NOT3 IN4 O9 AND4
XAND11 NOT1 IN2 NOT3 IN4 O10 AND4
XAND12 IN1 IN2 NOT3 IN4 O11 AND4
XAND13 NOT1 NOT2 IN3 IN4 O12 AND4
XAND14 IN1 NOT2 IN3 IN4 O13 AND4
XAND15 NOT1 IN2 IN3 IN4 O14 AND4
XAND16 IN1 IN2 IN3 IN4 O15 AND4


.ENDS DEC416

*---DFLIPFLOP--------------------------------------------------------------------------------

.SUBCKT DFLIPFLOP D Q


XNOT1 D NOTD NOT
XNOT2 CLK NOTCLK NOT

XNAND1 D NOTCLK NAND1 NAND
XNAND2 NOTCLK NOTD NAND2 NAND
XNAND3 NAND1 QNOT1 Q1 NAND
XNAND4 Q1 NAND2 QNOT1 NAND

XNAND5 Q1 CLK NAND5 NAND
XNAND6 CLK QNOT1 NAND6 NAND
XNAND7 NAND5 QNOT Q NAND
XNAND8 Q NAND6 QNOT NAND

.ENDS DFLIPFLOP

*---PC--------------------------------------------------------------------------------

.SUBCKT PC IN1 IN2 IN3 IN4 OUT1 OUT2 OUT3 OUT4


XFLIPFLOP0 IN1 OUT1 DFLIPFLOP
XFLIPFLOP1 IN2 OUT2 DFLIPFLOP
XFLIPFLOP2 IN3 OUT3 DFLIPFLOP
XFLIPFLOP3 IN4 OUT4 DFLIPFLOP


.ENDS PC


*---HA--------------------------------------------------------------------------------

.SUBCKT HA INA INB S COUT 

XXOR INA INB S XOR
XAND INA INB COUT AND


.ENDS HA

*---FA--------------------------------------------------------------------------------

.SUBCKT FA A B C S COUT

XHA1 A B S1 C1 HA
XHA2 S1 C S C2 HA

XOR C1 C2 COUT OR

.ENDS FA

*---ALU--------------------------------------------------------------------------------

.SUBCKT ALU Q0 Q1 Q2 Q3 D0 D1 D2 D3

VDD1 ADD1 0 1.1
XFA1 Q0 ADD1 0 D0 COUT1 FA
XFA2 Q1 COUT1 0 D1 COUT2 FA
XFA3 Q2 COUT2 0 D2 COUT3 FA
XFA4 Q3 COUT3 0 D3 COUT4 FA


.ENDS ALU


*------------------------------------------------------------------------------------

.END